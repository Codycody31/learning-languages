module main

fn main() {
	// the fuck can I not do camel case
	curse_words := ['shitty', 'fucking', 'smelly']
	for curse in curse_words {
		println('Hello ${curse} world!')
	}
}
